//******************************************************************************
//
//******************************************************************************


`include "PODES_M0A_reg_define.h"
`include "AMY_reg_define.h"


module testcase ();

//blank testcase. 
//simulation just runs test program from ROM.

endmodule
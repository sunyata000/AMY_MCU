//******************************************************************************
//
//******************************************************************************


`include "PODES_M0A_reg_define.h"
`include "AMY_reg_define.h"


module testcase (sim_done);

output sim_done;

reg sim_done = 1'b1;

endmodule
